module listiny_struct

pub struct SoundState {
pub mut:
	index      int
	is_playing bool
	is_paused  bool
}
