module listiny_button_fn

/*
import listiny_struct { App }

pub fn btn_page_back(mut app App, x voidptr) {
	after := app.form.page_index - 1
	if after == -1 {
		app.form.page_index = app.nb_page - 1
	} else {
		app.form.page_index = after
	}
}*/
