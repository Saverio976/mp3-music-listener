module yt_dl_button_fn

/*
import yt_dl_struct { App }

pub fn btn_page_next(mut app App, x voidptr) {
	after := app.form.page_index + 1
	if after == app.nb_page {
		app.form.page_index = 0
	} else {
		app.form.page_index = after
	}
}*/
